interface inter #(parameter N = 5) ();   // note: parameter list AFTER the name
    logic [N-1:0] a;
    logic [N-1:0] b;
    logic [N-1:0] out;
endinterface
