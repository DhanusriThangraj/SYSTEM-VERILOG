interface inter();
  logic clk;
  logic [2:0]addr;
  logic [3:0]data;
endinterface
