xcelium> run
TIME	CLK	RESET	J	K	Q	Qbar	
0	    0	x	x	x	x	x
5	    1	1	x	x	0	1
10	  0	0	x	x	0	1
15   	1	0	0	1	0	1
20  	0	0	0	0	0	1
25  	1	0	1	1	1	0
30	  0	0	1	0	1	0
Simulation complete via $finish(1) at time 31 NS + 0
./test.sv:22      #1;$finish;  
xcelium> exit
TOOL:	xrun	23.09-s001: Exiting on Sep 07, 2025 at 08:19:55 EDT  (total: 00:00:01)
Done
