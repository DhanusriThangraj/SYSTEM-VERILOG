Compiler version U-2023.03-SP2_Full64; Runtime version U-2023.03-SP2_Full64;  Sep  8 05:03 2025
A=x B=x SUM=x
A=10 B=15 SUM=25
           V C S   S i m u l a t i o n   R e p o r t 
Time: 0 ns
CPU Time:      0.400 seconds;       Data structure size:   0.0Mb
Mon Sep  8 05:04:00 2025
Done
