
module func;
  initial begin
    display();
  end
  
  function void  display();
      $display("DHANU");
    endfunction
endmodule

// output
Compiler version U-2023.03-SP2_Full64; Runtime version U-2023.03-SP2_Full64;  Sep 29 00:44 2025
DHANU
           V C S   S i m u l a t i o n   R e p o r t 
Time: 0 ns
CPU Time:      0.350 seconds;       Data structure size:   0.0Mb
Mon Sep 29 00:44:24 2025
Done
