module example;
  initial begin
    repeat(5)begin
      $display("GOOD MORNING");
      $display("------------");
    end
  end
endmodule
// output
Compiler version U-2023.03-SP2_Full64; Runtime version U-2023.03-SP2_Full64;  Aug 30 12:45 2025
GOOD MORNING
------------
GOOD MORNING
------------
GOOD MORNING
------------
GOOD MORNING
------------
GOOD MORNING
------------
           V C S   S i m u l a t i o n   R e p o r t 
Time: 0 ns
CPU Time:      0.420 seconds;       Data structure size:   0.0Mb
Sat Aug 30 12:45:35 2025
Done

