module byte_;
  byte a; 
  byte b;
  byte c;
  byte d;
  byte e;
  byte f;

  initial begin
    a ='bxxz;                 // sized
    $display("a = %b", a);

    b = 'bxxxxxzzzzx;
    $display("b = %b", b);

    c ='bxxzzz1x;  
    $display("c = %b", c);

    d ='bxxzz010x;     
    $display("d = %b", d);

    e = 'bxxzz100111;  
    $display("e = %b", e);

    f = 'bxxzz100110010;   
    $display("f = %b", f);
  end
endmodule

// output
xcelium> run
a = 00000000
b = 00000000
c = 00000010
d = 00000100
e = 00100111
f = 00110010
xmsim: *W,RNQUIE: Simulation is complete.
xcelium> exit
