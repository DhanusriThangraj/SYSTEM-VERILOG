# run -all
# DATA=12 ADDR=4
# DATA=14 ADDR=5
# ** Note: $finish    : testbench.sv(20)
