Compiler version U-2023.03-SP2_Full64; Runtime version U-2023.03-SP2_Full64;  Sep  7 08:28 2025
Time	A	B		OUT
0	110	11111		110	
10	11110	10011		10010	
$finish called from file "top.sv", line 15.
$finish at simulation time                   11
           V C S   S i m u l a t i o n   R e p o r t 
Time: 11 ns
CPU Time:      0.360 seconds;       Data structure size:   0.0Mb
Sun Sep  7 08:28:10 2025
Done
