xcelium> source /xcelium23.09/tools/xcelium/files/xmsimrc
xcelium> run
Time	A	sel	Y	
0	x	x	x	
1	1010	0	0	
13	1010	1	1	
28	1010	10	0	
48	1010	11	1	
Simulation complete via $finish(1) at time 49 NS + 0
./top.sv:15     #1;$finish;
xcelium> exit
TOOL:	xrun	23.09-s001: Exiting on Sep 07, 2025 at 08:27:05 EDT  (total: 00:00:01)
Done
