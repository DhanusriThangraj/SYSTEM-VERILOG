xcelium> source /xcelium23.09/tools/xcelium/files/xmsimrc
xcelium> run
A	B	C	SUM	SUB
x	x	x	x	 x
11	x	x	x	 x
11	1010	x	1101	 x
11	1010	10	1101	11
Simulation complete via $finish(1) at time 16 NS + 0
./testbench.sv:20     #1;$finish;
xcelium> exit
TOOL:	xrun	23.09-s001: Exiting on Sep 08, 2025 at 06:35:27 EDT  (total: 00:00:01)
Done
