interface inter;
  logic [3:0]a;
  logic [1:0]sel;
  logic y;
endinterface
